* C:\Users\satyam\Desktop\LT Spice\Nand.cir
*
.include C:\Users\satyam\Desktop\LT Spice\180nm_model.txt
vdd 1 0 dc 1.8
* pulse_source pulse(Voff Von Delay Rise_time fall_time On_time time_period Cycles)
vA 2 0 pulse(0 1.8 0n 0.1n 0.1n 2n 4n)
vB 3 0 pulse(0 1.8 1n 0.1n 0.1n 2n 4n)
* device_name Drain Gate source substrate Device_model channel_width channel Height

MP0 4 2 1 1 P_180 w=4u l=.18u
MP1 4 3 1 1 P_180 w=4u l=.18u

MN0 4 2 5 0 N_180 w=2u l=.18u
MN1 5 3 0 0 N_180 w=2u l=.18u

MP2 C 4 1 1 P_180 w=4u l=.18u
MN2 C 4 0 0 N_180 w=2u l=.18u


MP3 7 2 1 1 P_180 w=4u l=.18u
MP4 7 4 1 1 P_180 w=4u l=.18u

MN3 7 2 6 0 N_180 w=2u l=.18u
MN4 6 4 0 0 N_180 w=2u l=.18u


MP5 9 3 1 1 P_180 w=4u l=.18u
MP6 9 4 1 1 P_180 w=4u l=.18u

MN5 9 3 8 0 N_180 w=2u l=.18u
MN6 8 4 0 0 N_180 w=2u l=.18u


MP7 S 7 1 1 P_180 w=4u l=.18u
MP8 S 9 1 1 P_180 w=4u l=.18u

MN7 S 7 10 0 N_180 w=2u l=.18u
MN8 10 9 0 0 N_180 w=2u l=.18u

.tran 0 50n

** Delay of A to S
**Tphl
.meas tran tpra
+ TRIG V(2) VAL = '1.8/2' RISE = 1
+ TARG V(S) VAL = '1.8/2' FALL = 1
** Tplh
.meas tran tpfa
+ TRIG V(2) VAL = '1.8/2' FALL = 1
+ TARG V(S) VAL = '1.8/2' RISE = 1

.meas tran tpd_A_S param=(tpra+tpfa)/2


** Delay of S to B

.meas tran tprb
+ TRIG V(S) VAL = '1.8/2' FALL = 1
+ TARG V(3) VAL = '1.8/2' RISE = 1

.meas tran tpfb
+ TRIG V(S) VAL = '1.8/2' RISE = 1
+ TARG V(3) VAL = '1.8/2' FALL = 1

.meas tran tpd_S_B param=(tprb+tpfb)/2
