
* C:\Users\satyam\Desktop\LT Spice\Nand.cir
*
.include C:\Users\satyam\Desktop\LT Spice\180nm_model.txt
vdd 1 0 dc 1.8
* pulse_source pulse(Voff Von Delay Rise_time fall_time On_time time_period Cycles)
va 2 0 pulse(0 1.8 0n 0.1n 0.1n 10n 20n)
vb 3 0 pulse(0 1.8 2n 0.1n 0.1n 10n 20n)
vc 4 0 pulse(0 1.8 4n 0.1n 0.1n 10n 20n)
* device_name Drain Gate source substrate Device_model channel_width channel Height
MP0 Vout 2 1 1 P_180 w=20u l=.18u
MP1 Vout 3 1 1 P_180 w=20u l=.18u
MP2 Vout 4 1 1 P_180 w=20u l=.18u

MN0 Vout 2 6 0 N_180 w=5u l=.18u
MN1 6 3 5 0 N_180 w=5u l=.18u
MN2 5 4 0 0 N_180 w=5u l=.18u
.tran 0 100n
*.dc va 0 1.8
.print tran v(Vout) v(4) v(2) v(3)
