*
.include 180nm_model.txt
.param SUPPLY=1.8V
*X1
M1 3 2 1 1 P_180 w=0.72u l=.18u
M2 3 2 0 0 N_180 w=0.36u l=.18u
*X2
M3 4 3 1 1 P_180 w=2.880u l=.18u
M4 4 3 0 0 N_180 w=1.440u l=.18u
*X3 Same
M5 5 4 1 1 P_180 w=11.520u l=.18u
M6 5 4 0 0 N_180 w=5.760u l=.18u
*X4
M7 6 5 1 1 P_180 w=46.080u l=.18u
M8 6 5 0 0 N_180 w=23.040u l=.18u
*X5
M9 7 6 1 1 P_180 w=184.320u l=.18u
M10 7 6 0 0 N_180 w=92.160u l=.18u
*X6 Same
M11 8 4 1 1 P_180 w=11.520u l=.18u
M12 8 4 0 0 N_180 w=5.760u l=.18u
Cdelay 8 0 135.67859ff
Vdd 1 0 DC 1.8v
Vin 2 0 PULSE(0 1.8 0n 0.1n 0.1n 10n 20n)
.tran 0 100ns
*-----------------------------------------------------------
*** Delay Calculations ***
*-----------------------------------------------------------
***** 4 to 5 Delay------------------------------------------
*** rising prop delay
.measure tran tpdr45
+ TRIG v(4) VAL='SUPPLY/2' RISE=2
+ TARG v(5) VAL='SUPPLY/2' FALL=2
*** falling prop delay
.measure tran tpdf45
+ TRIG v(4) VAL='SUPPLY/2' FALL=2
+ TARG v(5) VAL='SUPPLY/2' RISE=2
.measure tran avg_tpd45_inps param=(tpdr45+tpdf45)/2p
*** average prop delay (in ps)
***** 4 to 8 Delay------------------------------------------
*** rising prop delay
.measure tran tpdr48
+ TRIG v(4) VAL='SUPPLY/2' RISE=2
+ TARG v(8) VAL='SUPPLY/2' FALL=2
*** falling prop delay
.measure tran tpdf48
+ TRIG v(4) VAL='SUPPLY/2' FALL=2
+ TARG v(8) VAL='SUPPLY/2' RISE=2
.measure tran avg_tpd48_inps param=(tpdr48+tpdf48)/2p
*** average prop delay (in ps)

.measure tran relation param=135.678/(46080+23040)
