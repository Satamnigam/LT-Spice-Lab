* C:\Users\satyam\Desktop\LT Spice\Nand.cir
* select_line >> v(4) V0>>v(3) V1>>v(2)
.include C:\Users\satyam\Desktop\LT Spice\180nm_model.txt
vdd 1 0 dc 1.8
* pulse_source pulse(Voff Von Delay Rise_time fall_time On_time time_period Cycles)
v1 2 0 pulse(0 1.8 0n 0.1n 0.1n 10n 20n)
v0 3 0 pulse(0 1.8 5n 0.1n 0.1n 10n 20n)
v2 4 0 pulse(0 1.8 6n 0.1n 0.1n 8n 20n)
* device_name Drain Gate source substrate Device_model channel_width channel Height

*First And gate
MP0 7 2 1 1 P_180 w=20u l=.18u
MP1 7 4 1 1 P_180 w=20u l=.18u
MP2 8 7 1 1 P_180 w=20u l=.18u

MN0 7 2 12 0 N_180 w=5u l=.18u
MN1 12 4 0 0 N_180 w=5u l=.18u
MN2 8 7 0 0 N_180 w=5u l=.18u

*not gate
MP3 11 4 1 1 P_180 w=20u l=.18u
MN3 11 4 0 0 N_180 w=5u l=.18u

*second and gate
MP4 5 11 1 1 P_180 w=20u l=.18u
MP5 5 3 1 1 P_180 w=20u l=.18u
MP6 9 5 1 1 P_180 w=20u l=.18u

MN4 5 11 4 0 N_180 w=5u l=.18u
MN5 4 3 0 0 N_180 w=5u l=.18u
MN6 9 5 0 0 N_180 w=5u l=.18u

*OR gate
MP7 6 8 1 1 P_180 w=20u l=.18u
MP8 10 9 6 6 P_180 w=20u l=.18u
MP9 Vout 10 1 1 P_180 w=20u l=.18u

MN7 10 8 0 0 N_180 w=5u l=.18u
MN8 10 9 0 0 N_180 w=5u l=.18u
MN9 Vout 10 0 0 N_180 w=5u l=.18u

.tran 0 100n

*.dc va 0 1.8
.print tran v(Vout) v(2) v(3) v(4)
.meas tran tar
+ TRIG V(2) VAL = '1.8/2' FALL = 1
+ TARG V(Vout) VAL = '1.8/2' RISE = 1
.meas tran taf
+ TRIG V(2) VAL = '1.8/2' RISE = 1
+ TARG V(Vout) VAL = '1.8/2' FALL = 1
.measure tran avg_tpda param=(tar+taf)/2p

.meas tran tprb
+ TRIG V(3) VAL = '1.8/2' FALL = 1
+ TARG V(Vout) VAL = '1.8/2' RISE = 1
.meas tran tpfb
+ TRIG V(3) VAL = '1.8/2' RISE = 1
+ TARG V(Vout) VAL = '1.8/2' FALL = 1
.measure tran avg_tpdb param=(tprb+tpfb)/2p
