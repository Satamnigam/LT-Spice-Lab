
* C:\Users\satyam\Desktop\LT Spice\Nand.cir
*
.include C:\Users\satyam\Desktop\LT Spice\180nm_model.txt
vdd 1 0 dc 1.8
* pulse_source pulse(Voff Von Delay Rise_time fall_time On_time time_period Cycles)
va A 0 pulse(0 1.8 0n 0.1n 0.1n 5n 20n)
vb B 0 pulse(0 1.8 3n 0.1n 0.1n 10n 20n)
vc S 0 pulse(0 1.8 7n 0.1n 0.1n 8n 20n)

* device_name Drain Gate source substrate Device_model channel_width channel Height
*STAGE 1
MP0 Sbar S 1 1 P_180 w=0.72u l=.18u
MP1 Sbar S 1 1 P_180 w=0.72u l=.18u
MN0 Sbar S 3 0 N_180 w=0.36u l=.18u
MN1 3 S 0 0 N_180 w=0.36u l=.18u

MP4 y B 1 1 P_180 w=0.72u l=.18u
MP5 y S 1 1 P_180 w=0.72u l=.18u
MN4 y B 5 0 N_180 w=0.72u l=.18u
MN5 5 S 0 0 N_180 w=0.72u l=.18u

*STAGE 2
MP2 x A 1 1 P_180 w=1.648u l=.18u
MP3 x Sbar 1 1 P_180 w=1.648u l=.18u
MN2 x A 4 0 N_180 w=0.824u l=.18u
MN3 4 Sbar 0 0 N_180 w=0.824u l=.18u

*STAGE 3
MP6 O x 1 1 P_180 w=3.774u l=.18u
MP7 O y 1 1 P_180 w=3.774u l=.18u
MN6 O x 6 0 N_180 w=1.887u l=.18u
MN7 6 y 0 0 N_180 w=1.887u l=.18u

.tran 0 100n
*.dc va 0 1.8
.print tran v(A) v(B) v(S) v(O)
.meas tran tar
+ TRIG V(A) VAL = '1.8/2' FALL = 1
+ TARG V(O) VAL = '1.8/2' RISE = 1
.meas tran taf
+ TRIG V(A) VAL = '1.8/2' RISE = 1
+ TARG V(O) VAL = '1.8/2' FALL = 1
.measure tran avg_tpda param=(tar+taf)/2p

.meas tran tprb
+ TRIG V(B) VAL = '1.8/2' FALL = 1
+ TARG V(O) VAL = '1.8/2' RISE = 1
.meas tran tpfb
+ TRIG V(B) VAL = '1.8/2' RISE = 1
+ TARG V(O) VAL = '1.8/2' FALL = 1
.measure tran avg_tpdb param=(tprb+tpfb)/2p
